module alu#(
	parameter DW = 32,
	parameter AW = 32
)(
	input	logic [3-1:0]	alu_sel,
	input	logic [DW-1:0]	op1,
	input	logic [DW-1:0]	op2,
	output 	logic [DW-1:0]	res // result
);

	always_comb begin
		case(alu_sel)
			3'b000: res  = 'h0;
			3'b001: res  = op1 + op2;

			default: res = 'h0;
		endcase
	end


endmodule
