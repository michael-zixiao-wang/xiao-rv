`define XIAO_RV 0321 // my birthday

`define RISC_ISA 32
`define	PC_RST_ADDR 32'h0000_0000

